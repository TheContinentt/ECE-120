-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION lab6_struct_config OF lab6 IS
   FOR struct
   END FOR;
END lab6_struct_config;
